

package shared_pkg;

class shared_pkg_c;
    static integer correct_count = 0;
    static integer error_count = 0;

    static bit test_finished;
endclass
endpackage